module pwm (
  input i_clk,
  input i_en,
  output reg o_pwm
);

  // Today's episode was amazing
endmodule